//TODO will tie everything the in the decode stage together