module jzjpcc_execute
#(
	parameter int PC_MAX_B
)
(
);

endmodule