module jzjpcc_mem_processor
(
	//Inputs
	//TODO needs funct3
	input logic [31:0] aluResult_execute,
	input logic [31:0] rs2_execute,
	
	//Outputs
	output logic [31:0] memDataToWrite_execute,
	output logic [3:0] memByteMask_execute
);

//TODO

endmodule