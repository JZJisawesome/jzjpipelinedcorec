module jzjpcc
(
	input logic clock,
	input logic reset,//Asynchronous
	
	output logic [31:0] register31Value//For testing
);
/* Connections */

/* Modules */
//Stages

//Common modules

endmodule