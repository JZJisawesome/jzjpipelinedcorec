interface jzjpcc_memory_if
();

endinterface